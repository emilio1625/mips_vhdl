library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

entity control_unit is
  port (
    clock
  );
end entity;

architecture arch of control_unit is

begin

end architecture;
